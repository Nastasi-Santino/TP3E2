module antiBounce (
    input clk,
    input rst,
    input wire rows[3:0],
    output reg validatedRows[3:0]
)




endmodule